class axi_environment extends uvm_env;

endclass
