interface axi_interface (
    input logic aclk,
    input logic arestn
);
endinterface
